module tenthirty(
    input clk,
    input rst_n, //negedge reset
    input btn_m, //bottom middle
    input btn_r, //bottom right
    output reg [7:0] seg7_sel,
    output reg [7:0] seg7,   //segment right
    output reg [7:0] seg7_l, //segment left
    output reg [2:0] led // led[0] : dealer win, led[1] : player win, led[2] : done
);

//================================================================
//   PARAMETER
//================================================================


//================================================================
//   d_clk
//================================================================
//frequency division
reg [24:0] counter; 
wire dis_clk; //seg display clk
wire d_clk  ; //division clk

//====== frequency division ======
always@(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        counter <= 0;
    end
    else begin
        counter <= counter + 1;
    end
end

//================================================================
//   REG/WIRE
//================================================================
//seg7_temp
reg [7:0] seg7_temp[0:7];

//================================================================
//   FLAG
//================================================================


//================================================================
//   FSM
//================================================================

//================================================================
//   I/O
//================================================================

reg  pip;
wire empty;
wire [3:0] number;

//================================================================
//   DESIGN
//================================================================




//================================================================
//   SEGMENT
//================================================================


//================================================================
//   LED
//================================================================

//================================================================
//   LUT
//================================================================
LUT inst_LUT (.clk(d_clk), .rst_n(rst_n), .pip(pip), .number(number), .empty(empty));

endmodule 